`timescale 1ns / 1ps
`include "constants.vh"
`include "helpers.vh"


module fadder_tb;

    reg [31:0] a, b, out;

    fadders UUT(.*);
    
    initial begin
        `TB_BEGIN;
        
        // -27.12 + 35.8 = 8.68
        a <= 32'b11000001110110001111010111000011;
        b <= 32'b01000010000011110011001100110011;
        #1 assert(out == 32'b01000001000010101110000101000110) else $error("[1]");
        
        // 0.005134 + 0.01954 = 0.24674
        a <= 32'b00111011101010000011101100011101;
        b <= 32'b00111100101000000001001001011010;
        #1 assert(out == 32'b00111100110010100010000100100001) else $error("[2]");
        
        // 0.4739 + 0.21005 = 0.68395
        a <= 32'b00111110111100101010001100000101;
        b <= 32'b00111110010101110001011101011001;
        #1 assert(out == 32'b00111111001011110001011101011000) else $error("[3]");
        
        // 0.08549374 + 0.09638762 = 0.18188136
        a <= 32'b00111101101011110001011101011000;
        b <= 32'b00111101110001010110011011011111;
        #1 assert(out == 32'b00111110001110100011111100011011) else $error("[4]");
        
        // 770059249123328 + 13.634336 = 770059249123345.634336 (770059249123328)
        a <= 32'b01011000001011110001011101011100;
        b <= 32'b01000001010110100010011000111110;
        #1 assert(out == 32'b01011000001011110001011101011100) else $error("[5]");
        
        // -429.613 + -982.119 = -1411.732
        a <= 32'b11000011110101101100111001110111;
        b <= 32'b11000100011101011000011110011110;
        #1 assert(out == 32'b11000100101100000111011101101100) else $error("[6]");
        
        `TB_END;
        $finish;
    end

endmodule
