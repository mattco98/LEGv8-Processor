`timescale 1ns / 1ps
`include "constants.vh"

module instruction_mem(

    );
endmodule
