`define FILE_BASE        "/home/matthew/Programming/LEGV8-Processor/LEGv8-Processor/instruction_sets/"
`define INSTRUCTION_FILE {`FILE_BASE, "general/instructions"}
`define RAM_FILE         {`FILE_BASE, "general/ram"}
`define REGISTERS_FILE   {`FILE_BASE, "general/registers"}

`define INSTRUCTION_FILE_DIVISION {`FILE_BASE, "division/division.instructions"}
`define RAM_FILE_DIVISION         {`FILE_BASE, "division/division.ram"}

`define INSTRUCTION_FILE_CMP {`FILE_BASE, "simple_compare/simple_compare.instructions"}
`define REGISTER_FILE_CMP    {`FILE_BASE, "simple_compare/simple_compare.registers"}