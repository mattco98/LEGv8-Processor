`define CYCLE 10