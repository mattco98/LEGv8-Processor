`define INSTRUCTION_FILE "C:\Users\matth\Documents\Programming\LEGV8-Processor\ARM-Processor\nonpipelined\sources\data\instructions"
`define RAM_FILE         "C:\Users\matth\Documents\Programming\LEGV8-Processor\ARM-Processor\nonpipelined\sources\data\ram"
`define REGISTERS_FILE   "C:\Users\matth\Documents\Programming\LEGV8-Processor\ARM-Processor\nonpipelined\sources\data\registers"