`define FILE_BASE        "/home/matthew/Programming/LEGV8-Processor/LEGv8-Processor/nonpipelined/sources/data/"
`define INSTRUCTION_FILE {`FILE_BASE, "instructions"}
`define RAM_FILE         {`FILE_BASE, "ram"}
`define REGISTERS_FILE   {`FILE_BASE, "registers"}

`define INSTRUCTION_MEM_TB_INSTR_FILE {`FILE_BASE, "instruction_mem_tb_instructions"}
`define REGISTER_MEM_TB_REGISTER_FILE {`FILE_BASE, "register_mem_tb_registers"}

`define INSTRUCTION_FILE_DIVISION {`FILE_BASE, "instructions_division"}
`define RAM_FILE_DIVISION         {`FILE_BASE, "ram_division"}