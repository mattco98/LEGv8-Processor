`define FILE_BASE        "C:/Users/matth/Documents/Programming/LEGV8-Processor/ARM-Processor/nonpipelined/sources/data/"
`define INSTRUCTION_FILE {`FILE_BASE, "instructions"}
`define RAM_FILE         {`FILE_BASE, "ram"}
`define REGISTERS_FILE   {`FILE_BASE, "registers"}

`define INSTRUCTION_MEM_TB_INSTR_FILE {`FILE_BASE, "instruction_mem_tb_instructions"}
`define REGISTER_MEM_TB_REGISTER_FILE {`FILE_BASE, "register_mem_tb_registers"}