`define FILE_BASE        "/home/matthew/Programming/LEGV8-Processor/LEGv8-Processor/instruction_sets/"
`define INSTRUCTION_FILE {`FILE_BASE, "general/instructions"}
`define RAM_FILE         {`FILE_BASE, "general/ram"}
`define REGISTERS_FILE   {`FILE_BASE, "general/registers"}

`define INSTRUCTION_FILE_DIVISION_UNSIGNED {`FILE_BASE, "division_unsigned/instructions"}
`define RAM_FILE_DIVISION_UNSIGNED         {`FILE_BASE, "division_unsigned/ram"}
`define REGISTER_FILE_DIVISION_UNSIGNED    {`FILE_BASE, "division_unsigned/registers"}

`define INSTRUCTION_FILE_DIVISION_SIGNED {`FILE_BASE, "division_signed/instructions"}
`define RAM_FILE_DIVISION_SIGNED         {`FILE_BASE, "division_signed/ram"}
`define REGISTER_FILE_DIVISION_SIGNED    {`FILE_BASE, "division_signed/registers"}

`define INSTRUCTION_FILE_CMP {`FILE_BASE, "simple_compare/instructions"}
`define REGISTER_FILE_CMP    {`FILE_BASE, "simple_compare/registers"}